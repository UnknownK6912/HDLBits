module top_module (
    input in,
    output out);

    wire mid;
    
    assign mid = in;
    assign out = mid;
    
endmodule
